module top_module(a,b,c,w,x,y,z);
    input wire a,b,c;
    output wire w,x,y,z;
    
    assign w=a;
    assign x=b;
    assign y=b;
    assign z=c;
    

endmodule