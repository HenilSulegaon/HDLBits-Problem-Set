module top_module ( input a, input b, output out );

    mod_a I1(a,b,out);
endmodule